module endScreen_rom (
	input logic clock,
	input logic [14:0] address,
	output logic [11:0] q
);

logic [11:0] memory [0:19199] /* synthesis ram_init_file = "./endScreen/endScreen.COE" */;

always_ff @ (posedge clock) begin
	q <= memory[address];
end

endmodule
